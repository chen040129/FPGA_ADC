// spi.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module spi (
		input  wire       clk_clk,                  //                                clk.clk
		input  wire       reset_reset_n,            //                              reset.reset_n
		input  wire       spislave_0_stsinkvalid,   //   spislave_0_avalon_streaming_sink.valid
		input  wire [7:0] spislave_0_stsinkdata,    //                                   .data
		output wire       spislave_0_stsinkready,   //                                   .ready
		input  wire       spislave_0_stsourceready, // spislave_0_avalon_streaming_source.ready
		output wire       spislave_0_stsourcevalid, //                                   .valid
		output wire [7:0] spislave_0_stsourcedata,  //                                   .data
		input  wire       spislave_0_mosi,          //                spislave_0_export_0.mosi
		input  wire       spislave_0_nss,           //                                   .nss
		inout  wire       spislave_0_miso,          //                                   .miso
		input  wire       spislave_0_sclk           //                                   .sclk
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> spislave_0:nreset

	SPIPhy #(
		.SYNC_DEPTH (2)
	) spislave_0 (
		.sysclk        (clk_clk),                         //              clock_sink.clk
		.nreset        (~rst_controller_reset_out_reset), //        clock_sink_reset.reset_n
		.mosi          (spislave_0_mosi),                 //                export_0.export
		.nss           (spislave_0_nss),                  //                        .export
		.miso          (spislave_0_miso),                 //                        .export
		.sclk          (spislave_0_sclk),                 //                        .export
		.stsourceready (spislave_0_stsourceready),        // avalon_streaming_source.ready
		.stsourcevalid (spislave_0_stsourcevalid),        //                        .valid
		.stsourcedata  (spislave_0_stsourcedata),         //                        .data
		.stsinkvalid   (spislave_0_stsinkvalid),          //   avalon_streaming_sink.valid
		.stsinkdata    (spislave_0_stsinkdata),           //                        .data
		.stsinkready   (spislave_0_stsinkready)           //                        .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
