library verilog;
use verilog.vl_types.all;
entity uart_tx_vlg_vec_tst is
end uart_tx_vlg_vec_tst;
