library verilog;
use verilog.vl_types.all;
entity clk_vlg_vec_tst is
end clk_vlg_vec_tst;
