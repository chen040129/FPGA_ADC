library verilog;
use verilog.vl_types.all;
entity uart_rx_vlg_vec_tst is
end uart_rx_vlg_vec_tst;
